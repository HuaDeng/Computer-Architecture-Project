/*CS 552 Project AND gate*/
module and_gate(in_1, in_2, out);
	
	input in_1, in_2;
	output out;

	and U(out, in_1, in_2);
endmodule 
